library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ECG_FPGA is
	port (
	);
end ECG_FPGA;

architecture RTL of ECG_FPGA is

begin

end architecture RTL;