library ieee;
use ieee.std_logic_1164.all;

package VGA_Char_Pkg is
	
	constant c_H_ACTIVE	: integer := 640;	--Horizontal screen width
	constant c_H_FP		: integer := 16;		--Horizontal front porch
	constant c_H_SP		: integer := 64;	--Horizontal sync width
	constant c_H_BP		: integer := 80;	--Horizontal back porch
	constant c_H_TOTAL	: integer := c_H_ACTIVE + c_H_FP + c_H_SP + c_H_BP;

	constant c_V_ACTIVE	: integer := 480;	--Vertical screen height
	constant c_V_FP		: integer := 3;		--Vertical front porch
	constant c_V_SP		: integer := 4;		--Vertical sync heigth
	constant c_V_BP		: integer := 13;		--Vertical back porch
	constant c_V_TOTAL	: integer := c_V_ACTIVE + c_V_FP + c_V_SP + c_V_BP;

	constant c_H_POL		: std_logic := '0';	--Horizontal sync polarity
	constant c_V_POL		: std_logic := '1';	--Vertical sync polarity
	constant c_BLANK_POL	: std_logic := '0';	--Blank polarity

	constant c_LIB_SIZE	: integer := 47;
	type t_CHAR is array(0 to 9) of std_logic_vector(0 to 7);
	type t_CHAR_ARRAY is array(0 to c_LIB_SIZE-1) of t_CHAR;

	constant c_LIB : t_CHAR_ARRAY := (
		0 => (	--char = '0'
			0 => "00000000",
			1 => "00111000",
			2 => "01001100",
			3 => "01010100",
			4 => "01100100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		1 => (	--char = '1'
			0 => "00000000",
			1 => "00010000",
			2 => "00110000",
			3 => "00010000",
			4 => "00010000",
			5 => "00010000",
			6 => "00010000",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		2 => (	--char = '2'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "00000100",
			4 => "00001000",
			5 => "00010000",
			6 => "00100000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),

		3 => (	--char = '3'
			0 => "00000000",
			1 => "01111100",
			2 => "00001000",
			3 => "00010000",
			4 => "00001000",
			5 => "00000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		4 => (	--char = '4'
			0 => "00000000",
			1 => "00001000",
			2 => "00011000",
			3 => "00101000",
			4 => "01001000",
			5 => "01111100",
			6 => "00001000",
			7 => "00001000",
			8 => "00000000",
			9 => "00000000"),

		5 => (	--char = '5'
			0 => "00000000",
			1 => "01111100",
			2 => "01000000",
			3 => "01111000",
			4 => "00000100",
			5 => "00000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		6 => (	--char = '6'
			0 => "00000000",
			1 => "00011000",
			2 => "00100000",
			3 => "01000000",
			4 => "01111000",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		7 => (	--char = '7'
			0 => "00000000",
			1 => "01111100",
			2 => "00000100",
			3 => "00001000",
			4 => "00010000",
			5 => "00100000",
			6 => "00100000",
			7 => "00100000",
			8 => "00000000",
			9 => "00000000"),

		8 => (	--char = '8'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "00111000",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		9 => (	--char = '9'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "00111100",
			5 => "00000100",
			6 => "00001000",
			7 => "00110000",
			8 => "00000000",
			9 => "00000000"),

		10 => (	--char = 'A'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01111100",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),

		11 => (	--char = 'B'
			0 => "00000000",
			1 => "01111000",
			2 => "01000100",
			3 => "01000100",
			4 => "01111000",
			5 => "01000100",
			6 => "01000100",
			7 => "01111000",
			8 => "00000000",
			9 => "00000000"),

		12 => (	--char = 'C'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000000",
			4 => "01000000",
			5 => "01000000",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		13 => (	--char = 'D'
			0 => "00000000",
			1 => "01110000",
			2 => "01001000",
			3 => "01000100",
			4 => "01000100",
			5 => "01000100",
			6 => "01001000",
			7 => "01110000",
			8 => "00000000",
			9 => "00000000"),	

		14 => (	--char = 'E'
			0 => "00000000",
			1 => "01111100",
			2 => "01000000",
			3 => "01000000",
			4 => "01111000",
			5 => "01000000",
			6 => "01000000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),

		15 => (	--char = 'F'
			0 => "00000000",
			1 => "01111100",
			2 => "01000000",
			3 => "01000000",
			4 => "01111000",
			5 => "01000000",
			6 => "01000000",
			7 => "01000000",
			8 => "00000000",
			9 => "00000000"),

		16 => (	--char = 'G'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000000",
			4 => "01011100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111100",
			8 => "00000000",
			9 => "00000000"),

		17 => (	--char = 'H'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "01111100",
			5 => "01000100",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),

		18 => (	--char = 'I'
			0 => "00000000",
			1 => "00111000",
			2 => "00010000",
			3 => "00010000",
			4 => "00010000",
			5 => "00010000",
			6 => "00010000",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		19 => (	--char = 'J'
			0 => "00000000",
			1 => "00011100",
			2 => "00001000",
			3 => "00001000",
			4 => "00001000",
			5 => "00001000",
			6 => "01001000",
			7 => "00110000",
			8 => "00000000",
			9 => "00000000"),

		20 => (	--char = 'K'
			0 => "00000000",
			1 => "01000100",
			2 => "01001000",
			3 => "01010000",
			4 => "01100000",
			5 => "01010000",
			6 => "01001000",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),

		21 => (	--char = 'L'
			0 => "00000000",
			1 => "01000000",
			2 => "01000000",
			3 => "01000000",
			4 => "01000000",
			5 => "01000000",
			6 => "01000000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),

		22 => (	--char = 'M'
			0 => "00000000",
			1 => "01000100",
			2 => "01101100",
			3 => "01010100",
			4 => "01010100",
			5 => "01000100",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),

		23 => (	--char = 'N'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01100100",
			4 => "01010100",
			5 => "01001100",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),

		24 => (	--char = 'O'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		25 => (	--char = 'P'
			0 => "00000000",
			1 => "01111000",
			2 => "01000100",
			3 => "01000100",
			4 => "01111000",
			5 => "01000000",
			6 => "01000000",
			7 => "01000000",
			8 => "00000000",
			9 => "00000000"),

		26 => (	--char = 'Q'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01010100",
			6 => "01001000",
			7 => "00110100",
			8 => "00000000",
			9 => "00000000"),

		27 => (	--char = 'R'
			0 => "00000000",
			1 => "01111100",
			2 => "01000100",
			3 => "01000100",
			4 => "01111000",
			5 => "01010000",
			6 => "01001000",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),

		28 => (	--char = 'S'
			0 => "00000000",
			1 => "00111100",
			2 => "01000000",
			3 => "01000000",
			4 => "00111000",
			5 => "00000100",
			6 => "00000100",
			7 => "01111000",
			8 => "00000000",
			9 => "00000000"),

		29 => (	--char = 'T'
			0 => "00000000",
			1 => "01111100",
			2 => "00010000",
			3 => "00010000",
			4 => "00010000",
			5 => "00010000",
			6 => "00010000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),

		30 => (	--char = 'U'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		31 => (	--char = 'V'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01000100",
			6 => "00101000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),

		32 => (	--char = 'W'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "01010100",
			5 => "01010100",
			6 => "01010100",
			7 => "00101000",
			8 => "00000000",
			9 => "00000000"),

		33 => (	--char = 'X'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "00101000",
			4 => "00010000",
			5 => "00101000",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),

		34 => (	--char = 'Y'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "00101000",
			5 => "00010000",
			6 => "00010000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),

		35 => (	--char = 'Z'
			0 => "00000000",
			1 => "01111100",
			2 => "00000100",
			3 => "00001000",
			4 => "00010000",
			5 => "00100000",
			6 => "01000000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),

		36 => (	--char = '?'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "00000100",
			4 => "00001000",
			5 => "00010000",
			6 => "00000000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),

		37 => (	--char = '='
			0 => "00000000",
			1 => "00000000",
			2 => "01111100",
			3 => "00000000",
			4 => "01111100",
			5 => "00000000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),

		38 => (	--char = '+'
			0 => "00000000",
			1 => "00010000",
			2 => "00010000",
			3 => "01111100",
			4 => "00010000",
			5 => "00010000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),

		39 => (	--char = '-'
			0 => "00000000",
			1 => "00000000",
			2 => "00000000",
			3 => "01111100",
			4 => "00000000",
			5 => "00000000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),

		40 => (	--char = '*'
			0 => "00000000",
			1 => "00000000",
			2 => "01010100",
			3 => "00111000",
			4 => "01111100",
			5 => "00111000",
			6 => "01010100",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),

		41 => (	--char = '/'
			0 => "00000000",
			1 => "00000000",
			2 => "00000100",
			3 => "00001000",
			4 => "00010000",
			5 => "00100000",
			6 => "01000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),

		42 => (	--char = '!'
			0 => "00000000",
			1 => "00010000",
			2 => "00010000",
			3 => "00010000",
			4 => "00010000",
			5 => "00000000",
			6 => "00000000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),

		43 => (	--char = 'Block'
			0 => "11111111",
			1 => "11111111",
			2 => "11111111",
			3 => "11111111",
			4 => "11111111",
			5 => "11111111",
			6 => "11111111",
			7 => "11111111",
			8 => "11111111",
			9 => "11111111"),

		44 => (	--char = 'Block Left'
			0 => "00000011",
			1 => "00000011",
			2 => "00000011",
			3 => "00000011",
			4 => "00000011",
			5 => "00000011",
			6 => "00000011",
			7 => "00000011",
			8 => "00000011",
			9 => "00000011"),

		45 => (	--char = 'Block Right'
			0 => "11000000",
			1 => "11000000",
			2 => "11000000",
			3 => "11000000",
			4 => "11000000",
			5 => "11000000",
			6 => "11000000",
			7 => "11000000",
			8 => "11000000",
			9 => "11000000"),

		46 => (	--char = ' '
			0 => "00000000",
			1 => "00000000",
			2 => "00000000",
			3 => "00000000",
			4 => "00000000",
			5 => "00000000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000")
	);

	type t_WR_REQ is record
		sel : integer range 0 to c_LIB_SIZE;
		scale : integer range 0 to 3;
		h_addr : integer range 0 to c_H_ACTIVE-1;
		v_addr : integer range 0 to c_V_ACTIVE-1;
	end record t_WR_REQ;

end package;